----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/02/2024 10:16:22 AM
-- Design Name: 
-- Module Name: MUX-4 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MUX_2_64bit is
    Port ( 
        clk             : in std_logic;
        s0              : in std_logic;
        a0, a1          : in std_logic_vector(31 downto 0);
        output          : out std_logic_vector(31 downto 0)
    );
end MUX_2_64bit;

architecture Behavioral of MUX_2_64bit is
begin
    process(clk, s0)
    begin
        if rising_edge(clk) then
            if s0 = '0' then
                output <= a0;
            elsif s0 = '1' then
                output <= a1;
            else output <= (others => '0');
            end if;
        end if;
    end process;
end Behavioral;
